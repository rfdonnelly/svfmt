function f(int a);
    return a * a;
endfunction

function g(int a, int b);
    return f(a, b) + b;
endfunction
